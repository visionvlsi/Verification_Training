module tb;

 reg [1:0]x;
 
 initial
  begin
   x=0;
    $display(x);
   
  
  end

 initial $display(x);
 initial $display(x);
 initial $display(x);
 initial $display(x);
 initial $display(x);
 
endmodule